`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:55 10/28/2022 
// Design Name: 
// Module Name:    control_path 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module control_path(
	input[5:0] opcode,
	input[5:0] funct,
	output reg[1:0] RDst,
	output reg[1:0] MReg,
	output reg[3:0] ALUOp,
	output reg RWrite,
	output reg MR,
	output reg MW,
	output reg ALUSr,
	output reg ALUSw,
	output reg Branch,
	output reg JAd,
	output reg JB
    );
	 always @(*)
		begin
			case(opcode)
			6'b000000:
				begin
					case(funct)
					6'b000000:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd1;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000001:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd1;
							ALUSw=1'b1;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					endcase
				end
			6'b000001:
				begin
					case(funct)
					6'b000000:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd2;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000001:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd3;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					endcase
				end
			6'b000010:
				begin
					case(funct)
					6'b000000:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b1;
							ALUOp=4'd4;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000001:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b1;
							ALUOp=4'd6;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000010:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd4;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000011:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd6;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000100:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b1;
							ALUOp=4'd7;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					6'b000101:
						begin
							RDst=2'd0;
							RWrite=1'b1;
							MR=1'b0;
							MW=1'b0;
							MReg=2'd0;
							ALUSr=1'b0;
							ALUOp=4'd7;
							ALUSw=1'b0;
							Branch=1'b0;
							JAd=1'b0;
							JB=1'b0;
						end
					endcase
				end
			6'b000011:
				begin
					RDst=2'd1;
					RWrite=1'b1;
					MR=1'b1;
					MW=1'b0;
					MReg=2'd1;
					ALUSr=1'b1;
					ALUOp=4'd8;
					ALUSw=1'b0;
					Branch=1'b0;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b000100:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b1;
					MReg=2'd0;
					ALUSr=1'b1;
					ALUOp=4'd8;
					ALUSw=1'b0;
					Branch=1'b0;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b000101:
				begin
					RDst=2'd0;
					RWrite=1'b1;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd9;
					ALUSw=1'b0;
					Branch=1'b0;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b000110:
				begin
					RDst=2'd0;
					RWrite=1'b1;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b1;
					ALUOp=4'd1;
					ALUSw=1'b0;
					Branch=1'b0;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b000111:
				begin
					RDst=2'd0;
					RWrite=1'b1;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b1;
					ALUOp=4'd1;
					ALUSw=1'b1;
					Branch=1'b0;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b001000:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b001001:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b1;
					JB=1'b0;
				end
			6'b001010:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b1;
				end
			6'b001011:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b1;
				end
			6'b001100:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b1;
				end
			6'b001101:
				begin
					RDst=2'd2;
					RWrite=1'b1;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd2;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b001110:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b0;
				end
			6'b001111:
				begin
					RDst=2'd0;
					RWrite=1'b0;
					MR=1'b0;
					MW=1'b0;
					MReg=2'd0;
					ALUSr=1'b0;
					ALUOp=4'd0;
					ALUSw=1'b0;
					Branch=1'b1;
					JAd=1'b0;
					JB=1'b0;
				end
			endcase
		end
endmodule

